<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-103.195,-1.57718,104.523,-109.993</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>-28,-57.5</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2</ID>
<type>AE_OR2</type>
<position>-27.5,-98</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_AND2</type>
<position>-34.5,-88</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>-20.5,-88</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>GA_LED</type>
<position>-42.5,-28</position>
<input>
<ID>N_in0</ID>60 </input>
<input>
<ID>N_in1</ID>9 </input>
<input>
<ID>N_in2</ID>6 </input>
<input>
<ID>N_in3</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>GA_LED</type>
<position>-32,-24</position>
<input>
<ID>N_in0</ID>59 </input>
<input>
<ID>N_in1</ID>7 </input>
<input>
<ID>N_in2</ID>8 </input>
<input>
<ID>N_in3</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AE_DFF_LOW_NT</type>
<position>-48,-41.5</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUTINV_0</ID>5 </output>
<output>
<ID>OUT_0</ID>6 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8</ID>
<type>BB_CLOCK</type>
<position>-68.5,-51</position>
<output>
<ID>CLK</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 500</lparam></gate>
<gate>
<ID>9</ID>
<type>AE_DFF_LOW_NT</type>
<position>-29.5,-46</position>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>7 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>10</ID>
<type>AI_XOR2</type>
<position>-35.5,-37</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_AND2</type>
<position>5.5,-12.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>GA_LED</type>
<position>-20.5,-18.5</position>
<input>
<ID>N_in0</ID>58 </input>
<input>
<ID>N_in1</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AE_DFF_LOW_NT</type>
<position>-8.5,-37</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>15 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>15</ID>
<type>AI_XOR2</type>
<position>10,-30</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AE_OR2</type>
<position>-5.5,-98.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>-13.5,-88.5</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_AND2</type>
<position>0.5,-88.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AI_XOR2</type>
<position>18.5,-30</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>-47.5,-27.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>-36,-23.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>-25,-18</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>-27.5,-54</position>
<gparam>LABEL_TEXT Controle</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AE_SMALL_INVERTER</type>
<position>-31,-82</position>
<input>
<ID>IN_0</ID>52 </input>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AE_SMALL_INVERTER</type>
<position>-35.5,-81</position>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>5.5,-7</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AE_SMALL_INVERTER</type>
<position>-1,-6</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>48</ID>
<type>AE_SMALL_INVERTER</type>
<position>-1,-8</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>50</ID>
<type>AE_SMALL_INVERTER</type>
<position>-3,-83</position>
<input>
<ID>IN_0</ID>52 </input>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>52</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-76,-19.5</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>59 </input>
<input>
<ID>IN_2</ID>58 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>-5,-3.5</position>
<gparam>LABEL_TEXT Calculo Decrescente</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>-6,-15</position>
<gparam>LABEL_TEXT Calculo Crescente</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>-27,-62</position>
<gparam>LABEL_TEXT Calculo Crescente</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>-37,-70.5</position>
<gparam>LABEL_TEXT Calculo Decrescente</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 90</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,-93,-20.5,-91</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>-93 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-26.5,-95,-26.5,-93</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-26.5,-93,-20.5,-93</points>
<intersection>-26.5 1</intersection>
<intersection>-20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-95,-28.5,-93</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-93 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-34.5,-93,-34.5,-91</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-34.5,-93,-28.5,-93</points>
<intersection>-34.5 1</intersection>
<intersection>-28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64.5,-51,-11.5,-51</points>
<connection>
<GID>8</GID>
<name>CLK</name></connection>
<intersection>-56 4</intersection>
<intersection>-32.5 3</intersection>
<intersection>-11.5 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-32.5,-51,-32.5,-47</points>
<connection>
<GID>9</GID>
<name>clock</name></connection>
<intersection>-51 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-56,-51,-56,-42.5</points>
<intersection>-51 1</intersection>
<intersection>-42.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-56,-42.5,-51,-42.5</points>
<connection>
<GID>7</GID>
<name>clock</name></connection>
<intersection>-56 4</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-11.5,-51,-11.5,-38</points>
<connection>
<GID>14</GID>
<name>clock</name></connection>
<intersection>-51 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,-42.5,-44,-34</points>
<intersection>-42.5 5</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-51,-34,-44,-34</points>
<intersection>-51 3</intersection>
<intersection>-44 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-51,-39.5,-51,-34</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-45,-42.5,-44,-42.5</points>
<connection>
<GID>7</GID>
<name>OUTINV_0</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-39.5,-42.5,-29</points>
<connection>
<GID>5</GID>
<name>N_in2</name></connection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45,-39.5,-42.5,-39.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25.5,-44,-25.5,-24</points>
<intersection>-44 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-31,-24,-25.5,-24</points>
<connection>
<GID>6</GID>
<name>N_in1</name></connection>
<intersection>-25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-26.5,-44,-25.5,-44</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>-25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34.5,-34,-34.5,-29.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-29.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-32,-29.5,-32,-25</points>
<connection>
<GID>6</GID>
<name>N_in2</name></connection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-34.5,-29.5,-32,-29.5</points>
<intersection>-34.5 0</intersection>
<intersection>-32 1</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-34,-36.5,-28</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-41.5,-28,-36.5,-28</points>
<connection>
<GID>5</GID>
<name>N_in1</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-27,-42.5,-6</points>
<connection>
<GID>5</GID>
<name>N_in3</name></connection>
<intersection>-11.5 1</intersection>
<intersection>-6 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-42.5,-11.5,2.5,-11.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>-42.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-42.5,-6,-3,-6</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>-42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32,-23,-32,-8</points>
<connection>
<GID>6</GID>
<name>N_in3</name></connection>
<intersection>-13.5 1</intersection>
<intersection>-8 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32,-13.5,2.5,-13.5</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>-32 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-32,-8,-3,-8</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>-32 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-79,-35.5,-40</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>-61.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-35.5,-61.5,-19.5,-61.5</points>
<intersection>-35.5 0</intersection>
<intersection>-19.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-19.5,-85,-19.5,-61.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-61.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-35,-3,-18.5</points>
<intersection>-35 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-19.5,-18.5,17.5,-18.5</points>
<connection>
<GID>13</GID>
<name>N_in1</name></connection>
<intersection>-3 0</intersection>
<intersection>9 18</intersection>
<intersection>17.5 20</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-5.5,-35,-3,-35</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-3 0</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>9,-27,9,-18.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>17.5,-27,17.5,-18.5</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-41.5,-101,-41.5,-44</points>
<intersection>-101 2</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-41.5,-44,-32.5,-44</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>-41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-41.5,-101,-27.5,-101</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>-41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-93.5,0.5,-91.5</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>-93.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-4.5,-95.5,-4.5,-93.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>-93.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-4.5,-93.5,0.5,-93.5</points>
<intersection>-4.5 1</intersection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6.5,-95.5,-6.5,-93.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>-93.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-13.5,-93.5,-13.5,-91.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>-93.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-13.5,-93.5,-6.5,-93.5</points>
<intersection>-13.5 1</intersection>
<intersection>-6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-27,11,-12.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-12.5,11,-12.5</points>
<connection>
<GID>11</GID>
<name>OUT</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-85,-33.5,-82</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33.5,-82,-33,-82</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-85,-35.5,-83</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1,-8,2.5,-8</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1,-6,2.5,-6</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-27,19.5,-7</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-7,19.5,-7</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18,-101.5,-18,-35</points>
<intersection>-101.5 2</intersection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-18,-35,-11.5,-35</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-18,-101.5,-5.5,-101.5</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>-18 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,-85.5,-0.5,-83</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1,-83,-0.5,-83</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>-0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-82,-28,-59.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>-82 1</intersection>
<intersection>-65.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29,-82,-21.5,-82</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>-28 0</intersection>
<intersection>-21.5 7</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-28,-65.5,-12.5,-65.5</points>
<intersection>-28 0</intersection>
<intersection>-12.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-12.5,-85.5,-12.5,-65.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-83 8</intersection>
<intersection>-65.5 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-21.5,-85,-21.5,-82</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-12.5,-83,-5,-83</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>-12.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-85.5,-14.5,-59</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>-59 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>10,-59,10,-33</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>-59 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-14.5,-59,10,-59</points>
<intersection>-14.5 0</intersection>
<intersection>10 1</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1.5,-85.5,1.5,-83</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-83 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>18.5,-83,18.5,-33</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>1.5,-83,18.5,-83</points>
<intersection>1.5 0</intersection>
<intersection>18.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-84,-14,-21.5,-14</points>
<intersection>-84 10</intersection>
<intersection>-21.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-21.5,-18.5,-21.5,-14</points>
<connection>
<GID>13</GID>
<name>N_in0</name></connection>
<intersection>-14 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-84,-18.5,-84,-14</points>
<intersection>-18.5 11</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-84,-18.5,-79,-18.5</points>
<connection>
<GID>52</GID>
<name>IN_2</name></connection>
<intersection>-84 10</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-90,-24,-33,-24</points>
<connection>
<GID>6</GID>
<name>N_in0</name></connection>
<intersection>-90 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-90,-24,-90,-19.5</points>
<intersection>-24 1</intersection>
<intersection>-19.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-90,-19.5,-79,-19.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>-90 3</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-83.5,-28,-43.5,-28</points>
<connection>
<GID>5</GID>
<name>N_in0</name></connection>
<intersection>-83.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-83.5,-28,-83.5,-20.5</points>
<intersection>-28 1</intersection>
<intersection>-20.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-83.5,-20.5,-79,-20.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-83.5 3</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,33.7192,492.369,-223.265</PageViewport></page 1>
<page 2>
<PageViewport>0,33.7192,492.369,-223.265</PageViewport></page 2>
<page 3>
<PageViewport>0,33.7192,492.369,-223.265</PageViewport></page 3>
<page 4>
<PageViewport>0,33.7192,492.369,-223.265</PageViewport></page 4>
<page 5>
<PageViewport>0,33.7192,492.369,-223.265</PageViewport></page 5>
<page 6>
<PageViewport>0,33.7192,492.369,-223.265</PageViewport></page 6>
<page 7>
<PageViewport>0,33.7192,492.369,-223.265</PageViewport></page 7>
<page 8>
<PageViewport>0,33.7192,492.369,-223.265</PageViewport></page 8>
<page 9>
<PageViewport>0,33.7192,492.369,-223.265</PageViewport></page 9></circuit>